//2 input and gate model
module and2(
    input a,
    input b,
    output y
);

assign y = a & b;
endmodule